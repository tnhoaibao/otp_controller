`timescale 1ns/10ps
module digtop (
	
);



memtop memtop_i (

);


endmodule